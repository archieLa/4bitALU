module display_output(in, display);

input [7:0] in;
output [7:0] display;

assign display = in;

endmodule 